** Profile: "SCHEMATIC1-test1"  [ C:\USERS\ZIM\DESKTOP\SMART CHARGER\Simulation\lm358 test-PSpiceFiles\SCHEMATIC1\test1.sim ] 

** Creating circuit file "test1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1.3ms 0 1us 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
